magic
tech sky130A
timestamp 1729095169
<< viali >>
rect 67 528 568 545
rect 66 18 567 35
<< metal1 >>
rect 61 545 574 548
rect 61 528 67 545
rect 568 528 574 545
rect 61 525 574 528
rect 85 271 90 297
rect 116 271 121 297
rect 141 274 313 295
rect 356 274 528 295
rect 548 271 553 297
rect 579 271 584 297
rect 60 35 573 38
rect 60 18 66 35
rect 567 18 573 35
rect 60 15 573 18
<< via1 >>
rect 90 271 116 297
rect 553 271 579 297
<< metal2 >>
rect 90 297 116 302
rect 553 297 579 302
rect 116 271 553 297
rect 90 266 116 271
rect 553 266 579 271
use inv  inv_0
timestamp 1729094408
transform 1 0 -156 0 1 -301
box 156 301 368 864
use inv  inv_1
timestamp 1729094408
transform 1 0 55 0 1 -301
box 156 301 368 864
use inv  inv_2
timestamp 1729094408
transform 1 0 266 0 1 -301
box 156 301 368 864
<< labels >>
flabel viali 187 531 187 531 0 FreeSans 160 0 0 0 vdd
port 0 nsew
flabel viali 184 23 184 23 0 FreeSans 160 0 0 0 gnd
port 1 nsew
flabel metal2 197 281 197 281 0 FreeSans 160 0 0 0 out
port 2 nsew
<< end >>
