** sch_path: /home/dwi/untitled.sch
**.subckt untitled
x1 net1 out GND ringosc3
V1 net1 GND 1.8
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/dwi/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/dwi/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/dwi/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/dwi/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.option wnflag=0
.option savecurrents
.control
save all
tran 1ps 10ns
plot out
op
.endc


**** end user architecture code
**.ends

* expanding   symbol:  ringosc3.sym # of pins=3
** sym_path: /home/dwi/ringosc3.sym
** sch_path: /home/dwi/ringosc3.sch
.subckt ringosc3 vdd out gnd
*.iopin vdd
*.iopin gnd
*.opin out
x1 vdd net1 net2 gnd inverterspice
x2 vdd net2 out gnd inverterspice
x3 vdd out net1 gnd inverterspice
.ends


* expanding   symbol:  inverterspice.sym # of pins=4
** sym_path: /home/dwi/.xschem/inverterspice.sym
** sch_path: /home/dwi/.xschem/inverterspice.sch
.subckt inverterspice vdd in out gnd
*.ipin in
*.opin out
*.ipin vdd
*.ipin gnd
XM2 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
